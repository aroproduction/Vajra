module main
// Main entry point

fn main() {
	println("Vajra 2.0 by GitHub Copilot")
	uci_loop()
}
