module main

import src

// Main entry point
fn main() {
	println("Vajra 2.0 by the Vajra Team")
	src.uci_loop()
}
